* D:\IV Semester\EW-2\Project-2\Audio_Amplifier.asc
.include "bc547.txt"

Q1 N004 N005 N006 0 BC547B
Q2 N002 0 N006 0 BC547B
R1 N001 N004 3k
R2 N001 N002 3k
R3 N006 N007 2k
V1 N001 0 12
V2 0 N007 12
V3 N005 0 SINE(0 10m 5k)
C1 N003 N002 100µ
* Q3 NC_01 NC_02 NC_03 0 TIP31C
* Q4 NC_04 NC_05 NC_06 0 TIP32C
.model NPN NPN
.model PNP PNP
* .lib C:\Users\jkoun\OneDrive\Documents\LTspiceXVII\lib\cmp\standard.bjt
.tran 20m
meas tran rptp pp v(N003) from=0 to =20m
.step temp 0 80 5
* .include "TIP31C.txt"
* .include "TIP32C.txt"
.backanno
.end